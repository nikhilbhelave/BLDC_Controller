`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:02:48 10/01/2016 
// Design Name: 
// Module Name:    pwm_nbv2 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pwm_nbv2(
    input [3:0] Q,
    input [3:0] D,
	 input clock ,
    output p
    );
	 wire [3:0] Q;
	 wire [3:0] D;
	 wire clock;
	 reg p;
	 for(
	 always @ (posedge clock)
	 Q <=


endmodule
